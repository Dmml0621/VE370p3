`timescale 1ns / 1ps

module Main_Memory_WB(
Address, WT, write, RD
    );

    input           write;
    input   [9:0]   Address;
    input   [127:0] WT;
    output  [127:0] RD;

    reg     [31:0] Memory[0:255];
    

    initial begin
        Memory[0] = 32'b11001000001111111010100100100110;
        Memory[1] = 32'b11001000001111111010100100100110;
        Memory[2] = 32'b10010001101100111101111110001001;
        Memory[3] = 32'b00011101101110011110000001110110;
        Memory[4] = 32'b11101010001100011010011110111001;
        Memory[5] = 32'b01110011000110011101101101010111;
        Memory[6] = 32'b01110100000101011010110010001000;
        Memory[7] = 32'b10101000100101011100011000100111;
        Memory[8] = 32'b00111111110111011101000111101110;
        Memory[9] = 32'b01100110010100101010111000000000;
        Memory[10] = 32'b11001000010110101100101011011111;
        Memory[11] = 32'b00011101010100101001010101110000;
        Memory[12] = 32'b10000010110111101010001110111111;
        Memory[13] = 32'b10000011110101101100110001000001;
        Memory[14] = 32'b01011111010111100011101110101110;
        Memory[15] = 32'b11001000011110000110010101101001;
        Memory[16] = 32'b00100101111100000000000011010110;
        Memory[17] = 32'b00111110111110000011111000011000;
        Memory[18] = 32'b10101010111101000100100111110111;
        Memory[19] = 32'b01100101011111000000011000101000;
        Memory[20] = 32'b11110100011101010111000010000110;
        Memory[21] = 32'b10101010111110110100111101001001;
        Memory[22] = 32'b00001111111000110000101110110110;
        Memory[23] = 32'b10010010101000110111000001011101;
        Memory[24] = 32'b01001001001011110000011110010011;
        Memory[25] = 32'b01011101001001110110100100101100;
        Memory[26] = 32'b10010010100011110111111011100001;
        Memory[27] = 32'b00000111100000010000100000001110;
        Memory[28] = 32'b00111100100010010110010111000000;
        Memory[29] = 32'b11111000000000010011001101111111;
        Memory[30] = 32'b01100111000011010000110010110000;
        Memory[31] = 32'b10111110100011000110101101011111;
        Memory[32] = 32'b10111000100001000001010110000001;
        Memory[33] = 32'b00000101000010000100000001101110;
        Memory[34] = 32'b11010000000000100110111011000001;
        Memory[35] = 32'b01011011000010100001100100011110;
        Memory[36] = 32'b00001111100001100100011011110000;
        Memory[37] = 32'b10010000101011100010000000111111;
        Memory[38] = 32'b00011101011001100101111111000000;
        Memory[39] = 32'b11101110011000100110111111001011;
        Memory[40] = 32'b11110010011010000010000000100101;
        Memory[41] = 32'b00100101111000000101011111110010;
        Memory[42] = 32'b10101100111011010010100100011101;
        Memory[43] = 32'b11111000011001010001111010010010;
        Memory[44] = 32'b01100111011111010101000001101110;
        Memory[45] = 32'b11001010011100010010010110000001;
        Memory[46] = 32'b00011001111110110101101001001110;
        Memory[47] = 32'b00000101110110110001110010100001;
        Memory[48] = 32'b11000010010101110010001100111111;
        Memory[49] = 32'b01011111010111110101010111010000;
        Memory[50] = 32'b11000100010101110011101000011111;
        Memory[51] = 32'b10100000110111110110111111100000;
        Memory[52] = 32'b00111111100100010101000101101110;
        Memory[53] = 32'b11101010000110000011011010000001;
        Memory[54] = 32'b01100010000100000110100001011010;
        Memory[55] = 32'b01110101100101000001101110110101;
        Memory[56] = 32'b10101000100111000111010001011011;
        Memory[57] = 32'b00000011100101000100000011000100;
        Memory[58] = 32'b01010111001110100001111100101011;
        Memory[59] = 32'b11001000001100100111100111100100;
        Memory[60] = 32'b01011101101110100000011000011010;
        Memory[61] = 32'b10010111101101100001000110010101;
        Memory[62] = 32'b10000010101111100111110101111000;
        Memory[63] = 32'b01111101001111100000101010100110;
        Memory[64] = 32'b11110000001100010111010001001001;
        Memory[65] = 32'b01100000101010010011001110100110;
        Memory[66] = 32'b00111111101000010000110000101001;
        Memory[67] = 32'b10111010111011010111101011010111;
        Memory[68] = 32'b01000001011001010011011100010000;
        Memory[69] = 32'b11010101010011010100000111111011;
        Memory[70] = 32'b10011010110000010111111001100100;
        Memory[71] = 32'b00000111110010110001110110001010;
        Memory[72] = 32'b10010101110010110100001101000101;
        Memory[73] = 32'b11011000010001110011010010111010;
        Memory[74] = 32'b01101101010011110101100001110101;
        Memory[75] = 32'b10110010110001100110111111011011;
        Memory[76] = 32'b00100010110010100011000000100100;
        Memory[77] = 32'b00101101010000000101011001101011;
        Memory[78] = 32'b11110000010010000010100110000100;
        Memory[79] = 32'b01100011011001000011111101011010;
        Memory[80] = 32'b10001111111001000101001011110101;
        Memory[81] = 32'b10011000111011000010010100111000;
        Memory[82] = 32'b00000101001000000101101111000111;
        Memory[83] = 32'b11000111001010100001110000001001;
        Memory[84] = 32'b01011010001000100010001010100110;
        Memory[85] = 32'b00000111101011100101011101101101;
        Memory[86] = 32'b10100000101101110001100010010010;
        Memory[87] = 32'b00111000001111110110101001111100;
        Memory[88] = 32'b11101111001110110101010110110011;
        Memory[89] = 32'b11100010001100010011001100001100;
        Memory[90] = 32'b00110101100110010110110011000011;
        Memory[91] = 32'b10101101100101010001100100101101;
        Memory[92] = 32'b10010010000111010111011111110010;
        Memory[93] = 32'b01010111000101010110000001011101;
        Memory[94] = 32'b11001111100110010001111010010010;
        Memory[95] = 32'b00011000100100110111100101100100;
        Memory[96] = 32'b00010101100100110000011110001011;
        Memory[97] = 32'b10001010010110100001001001000100;
        Memory[98] = 32'b01111010010101100111110111111011;
        Memory[99] = 32'b11110101110111100000101100110111;
        Memory[100] = 32'b10100000110101100111010011011100;
        Memory[101] = 32'b00111110111110000011001000000011;
        Memory[102] = 32'b11111111011100000000110110101100;
        Memory[103] = 32'b01000000011110000111110001100010;
        Memory[104] = 32'b01011101111111000011001010001101;
        Memory[105] = 32'b10011101111101000100010101010010;
        Memory[106] = 32'b00000010111111000111101110111100;
        Memory[107] = 32'b01010111011100100001110000010011;
        Memory[108] = 32'b11011000011010110100001111001100;
        Memory[109] = 32'b01101000111000110011011100100011;
        Memory[110] = 32'b10110111111011110001100011101101;
        Memory[111] = 32'b10101010100001110100111000010010;
        Memory[112] = 32'b01101100000001110011000110011101;
        Memory[113] = 32'b11110101000010110101011001110010;
        Memory[114] = 32'b01100010100000010010101010101100;
        Memory[115] = 32'b00001111100010010011110101000111;
        Memory[116] = 32'b10011111000001010101001101001000;
        Memory[117] = 32'b01000000000011010010010010110101;
        Memory[118] = 32'b11001101000001010111101101011011;
        Memory[119] = 32'b11011010100010000101100110010100;
        Memory[120] = 32'b00000010100010100010010001101011;
        Memory[121] = 32'b10100101000000100101001011100100;
        Memory[122] = 32'b11111000001011100001110100000010;
        Memory[123] = 32'b01101110001001100110101011001101;
        Memory[124] = 32'b11100111101011100101010000110010;
        Memory[125] = 32'b00111010101000100011001110111101;
        Memory[126] = 32'b00101101011010000110011101010011;
        Memory[127] = 32'b11010001011000000001100010001100;
        Memory[128] = 32'b01010010011001000011111101100011;
        Memory[129] = 32'b11001111111111000110000110001100;
        Memory[130] = 32'b10011000111101010001011000010110;
        Memory[131] = 32'b00010000011110010111100011111001;
        Memory[132] = 32'b11001111011100110000110100110110;
        Memory[133] = 32'b01111010010110110001001011001001;
        Memory[134] = 32'b00110100110101110111010001000111;
        Memory[135] = 32'b10100101110111110000111110101010;
        Memory[136] = 32'b00111000010111110101100101110101;
        Memory[137] = 32'b01111111010100110110010010011010;
        Memory[138] = 32'b11000011110110010000001101110100;
        Memory[139] = 32'b00011000110100010111110111101011;
        Memory[140] = 32'b10011101110111010010101000000100;
        Memory[141] = 32'b10000011000101000100010011001011;
        Memory[142] = 32'b01010010000111000111001100100101;
        Memory[143] = 32'b11001101101101000010111010111010;
        Memory[144] = 32'b00100000101100100100100001010101;
        Memory[145] = 32'b00110100101110100011011110011010;
        Memory[146] = 32'b10101111001100100000000101100000;
        Memory[147] = 32'b01101010001111100100111010101111;
        Memory[148] = 32'b11110101101101100011100100001000;
        Memory[149] = 32'b10100001101111100100010111110110;
        Memory[150] = 32'b00001010101100100000001000111001;
        Memory[151] = 32'b10010111001010000011110011010110;
        Memory[152] = 32'b01000001001010010100111100001001;
        Memory[153] = 32'b01001100101001010010000010100101;
        Memory[154] = 32'b10011111100011010111011011101010;
        Memory[155] = 32'b00000010100001010100101100010101;
        Memory[156] = 32'b00100110010010010010110111011010;
        Memory[157] = 32'b11111101010000110101001001110100;
        Memory[158] = 32'b01100000110010110000010110101011;
        Memory[159] = 32'b10100111110001111110101101000100;
        Memory[160] = 32'b10111011010001111101110010101011;
        Memory[161] = 32'b00101000010011111000000001100001;
        Memory[162] = 32'b11010101010000111110011111011110;
        Memory[163] = 32'b01010011110010001001100000010001;
        Memory[164] = 32'b00001110110000001010111011111110;
        Memory[165] = 32'b10010101011011001110000100100000;
        Memory[166] = 32'b01010000011001001001010110001111;
        Memory[167] = 32'b11001100011011001110101001000000;
        Memory[168] = 32'b11111111111010001010100010111111;
        Memory[169] = 32'b00110010111000101001011101010001;
        Memory[170] = 32'b10100101001010101110000010011110;
        Memory[171] = 32'b11111001001001101000111000100011;
        Memory[172] = 32'b01110010001111101101101111101100;
        Memory[173] = 32'b11000111101101101110010100000010;
        Memory[174] = 32'b00011001101110111000001011011101;
        Memory[175] = 32'b00011100000100011101110101111010;
        Memory[176] = 32'b11000101000100011010101110110001;
        Memory[177] = 32'b01010010100111011000010001001111;
        Memory[178] = 32'b11001110100101011111000010000000;
        Memory[179] = 32'b10100101100111011010111101101111;
        Memory[180] = 32'b00110000000100011100100011000000;
        Memory[181] = 32'b11101110000110111011011000011110;
        Memory[182] = 32'b01101011100100111000000111110001;
        Memory[183] = 32'b01110000100111111100111100111110;
        Memory[184] = 32'b10100101100111111011111011000001;
        Memory[185] = 32'b00001011010101101100000101001111;
        Memory[186] = 32'b01010110011110101100011110100000;
        Memory[187] = 32'b11000111111100101011100001111111;
        Memory[188] = 32'b01001000111110001100111010010001;
        Memory[189] = 32'b10011100111100001010001100011100;
        Memory[190] = 32'b10000011011111001111010011100011;
        Memory[191] = 32'b01101010011101001100101000001100;
        Memory[192] = 32'b11111100111101001010110111000110;
        Memory[193] = 32'b01100001111110001111001110111001;
        Memory[194] = 32'b00110010111000101000010000110110;
        Memory[195] = 32'b10111111011010101010100111011001;
        Memory[196] = 32'b01101011010001111101111100000111;
        Memory[197] = 32'b11010100110011111000000011101000;
        Memory[198] = 32'b10011101110001111110011001100111;
        Memory[199] = 32'b00001010010010111001100110001000;
        Memory[200] = 32'b10010110000010011000101001010110;
        Memory[201] = 32'b11010001000000011110011010111001;
        Memory[202] = 32'b01001000100011011001000101011110;
        Memory[203] = 32'b10111110100001011110111111000001;
        Memory[204] = 32'b00110011000011011110100000101111;
        Memory[205] = 32'b00101000000000011001011111100000;
        Memory[206] = 32'b11111101000010111110000100011111;
        Memory[207] = 32'b01110001101000101010110010010110;
        Memory[208] = 32'b10000110101001101101101001111000;
        Memory[209] = 32'b10011111001011101110010110100111;
        Memory[210] = 32'b00011000001001101000001001001000;
        Memory[211] = 32'b11000100001010101101110010100111;
        Memory[212] = 32'b01011011101000001010101100111001;
        Memory[213] = 32'b00001010101010001000011111010110;
        Memory[214] = 32'b10100100001001001111000000011001;
        Memory[215] = 32'b00110001011111001010111111100110;
        Memory[216] = 32'b11101010011111001100110100101000;
        Memory[217] = 32'b11101111111100001011001010000111;
        Memory[218] = 32'b00110011110110111010011001001000;
        Memory[219] = 32'b10101100010100111100100110110111;
        Memory[220] = 32'b10001101010111111011111001111001;
        Memory[221] = 32'b01010011110101111100000011010110;
        Memory[222] = 32'b11000110110111111100011100101101;
        Memory[223] = 32'b00001001110100111011100111100010;
        Memory[224] = 32'b00011000010100011100110000001100;
        Memory[225] = 32'b10000110010110011000101111010001;
        Memory[226] = 32'b01101011110101011111010101111110;
        Memory[227] = 32'b11111110110111011100001010110001;
        Memory[228] = 32'b10100101111101011010110001001111;
        Memory[229] = 32'b00110001011110001111101110001000;
        Memory[230] = 32'b11111110001100001000011000100111;
        Memory[231] = 32'b01101111101110101011000001111001;
        Memory[232] = 32'b01010001101111101111101110010110;
        Memory[233] = 32'b10011100101101101000110101111001;
        Memory[234] = 32'b00001011001111101111001010100110;
        Memory[235] = 32'b01010010001101101001010100001000;
        Memory[236] = 32'b11010100101010101000100111000111;
        Memory[237] = 32'b01001001101000001111111000101000;
        Memory[238] = 32'b10110100001010001001000011110011;
        Memory[239] = 32'b10110111000001001110011101011101;
        Memory[240] = 32'b01101011000001011111100110010010;
        Memory[241] = 32'b11111100100011011001110001101101;
        Memory[242] = 32'b01110101100000011110001110000010;
        Memory[243] = 32'b00000011000010111011010101001110;
        Memory[244] = 32'b10011110010000111101101011110001;
        Memory[245] = 32'b01000001010011111110110000111110;
        Memory[246] = 32'b11000000110001111001001111010001;
        Memory[247] = 32'b11011100110011111101011000001111;
        Memory[248] = 32'b00001011010000111010110010100000;
        Memory[249] = 32'b10100110010000011001101101101111;
        Memory[250] = 32'b11110101011010011101010110010000;
        Memory[251] = 32'b01101001111001001010001001011110;
        Memory[252] = 32'b11100110111011001101110110110001;
        Memory[253] = 32'b00110111011001001111100100001010;
        Memory[254] = 32'b00101001011010001010011011000101;
        Memory[255] = 32'b11001100011000101101000000100011;

    end

    assign RD = {Memory[{Address[9:4],2'b00}],Memory[{Address[9:4],2'b01}],Memory[{Address[9:4],2'b10}],Memory[{Address[9:4],2'b11}]};
    always @(Address, WT, write) begin
        if (write) begin
            Memory[{Address[9:4],2'b11}] = WT[31:0];
            Memory[{Address[9:4],2'b10}] = WT[63:32];
            Memory[{Address[9:4],2'b01}] = WT[95:64];
            Memory[{Address[9:4],2'b00}] = WT[127:96];
        end
    end

endmodule